LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY mux3 IS 
GENERIC(bits:INTEGER:=4);
PORT(
    in1,in2,in3,in4,in5,in6,in7,in8:IN STD_LOGIC_VECTOR(bits-1 DOWNTO 0);
    cin:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    out1:OUT STD_LOGIC_VECTOR(bits-1 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE arch OF mux3 IS 
begin
    out1<=in1 WHEN cin="000" ELSE in2 WHEN cin="001" ELSE in3 WHEN cin="010" ELSE in4 WHEN cin="011" ELSE in5 WHEN cin="100" ELSE in6 WHEN cin="101" ELSE in7 WHEN cin="110" ELSE in8 WHEN cin="111" ELSE in1;
END ARCHITECTURE;